library verilog;
use verilog.vl_types.all;
entity \register\ is
    port(
        \out\           : out    vl_logic_vector(9 downto 0);
        clk             : in     vl_logic
    );
end \register\;
