library verilog;
use verilog.vl_types.all;
entity tbb2 is
end tbb2;
