library verilog;
use verilog.vl_types.all;
entity shiba_vlg_vec_tst is
end shiba_vlg_vec_tst;
