library verilog;
use verilog.vl_types.all;
entity IMEM_vlg_vec_tst is
end IMEM_vlg_vec_tst;
