library verilog;
use verilog.vl_types.all;
entity alltb is
end alltb;
