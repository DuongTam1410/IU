library verilog;
use verilog.vl_types.all;
entity converterRGB_vlg_vec_tst is
end converterRGB_vlg_vec_tst;
