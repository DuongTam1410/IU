library verilog;
use verilog.vl_types.all;
entity tbb5 is
end tbb5;
