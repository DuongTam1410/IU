library verilog;
use verilog.vl_types.all;
entity all_vlg_vec_tst is
end all_vlg_vec_tst;
